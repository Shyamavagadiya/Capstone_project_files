library verilog;
use verilog.vl_types.all;
entity spi_testbench is
end spi_testbench;
