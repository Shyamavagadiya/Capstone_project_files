library verilog;
use verilog.vl_types.all;
entity spi_slave_test is
end spi_slave_test;
