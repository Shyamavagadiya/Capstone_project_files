library verilog;
use verilog.vl_types.all;
entity spi_master_test is
end spi_master_test;
